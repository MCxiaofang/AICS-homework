library verilog;
use verilog.vl_types.all;
entity tb_top_2 is
end tb_top_2;
